module ShiftRows(data_in, data_out);
    input [127:0] data_in;
    output [127:0] data_out;

    
endmodule