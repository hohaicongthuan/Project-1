module Second_Column_Mul(data_in, data_out);
    input [31:0] data_in;
    output [7:0] data_out;

    
endmodule